----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 10/15/2015 04:30:29 PM
-- Design Name: 
-- Module Name: invMixColumn - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

-- x9, x11, x13, x14 are the Gallois Multiplication Lookup Tables
-- Source: https://en.wikipedia.org/wiki/Rijndael_mix_columns#Galois_Multiplication_lookup_tables
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity x9 is
    Port ( byteIn : in STD_LOGIC_VECTOR(7 downto 0);
           byteOut : out STD_LOGIC_VECTOR(7 downto 0));
end x9;

architecture Behavioral of x9 is
begin
    process(byteIn)
    begin
        case byteIn is
            when x"00" => byteOut <= x"00";
            when x"01" => byteOut <= x"09";
            when x"02" => byteOut <= x"12";
            when x"03" => byteOut <= x"1B";
            when x"04" => byteOut <= x"24";
            when x"05" => byteOut <= x"2D";
            when x"06" => byteOut <= x"36";
            when x"07" => byteOut <= x"3F";
            when x"08" => byteOut <= x"48";
            when x"09" => byteOut <= x"41";
            when x"0A" => byteOut <= x"5A";
            when x"0B" => byteOut <= x"53";
            when x"0C" => byteOut <= x"6C";
            when x"0D" => byteOut <= x"65";
            when x"0E" => byteOut <= x"7E";
            when x"0F" => byteOut <= x"77";
            when x"10" => byteOut <= x"90";
            when x"11" => byteOut <= x"99";
            when x"12" => byteOut <= x"82";
            when x"13" => byteOut <= x"8B";
            when x"14" => byteOut <= x"B4";
            when x"15" => byteOut <= x"BD";
            when x"16" => byteOut <= x"A6";
            when x"17" => byteOut <= x"AF";
            when x"18" => byteOut <= x"D8";
            when x"19" => byteOut <= x"D1";
            when x"1A" => byteOut <= x"CA";
            when x"1B" => byteOut <= x"C3";
            when x"1C" => byteOut <= x"FC";
            when x"1D" => byteOut <= x"F5";
            when x"1E" => byteOut <= x"EE";
            when x"1F" => byteOut <= x"E7";
            when x"20" => byteOut <= x"3B";
            when x"21" => byteOut <= x"32";
            when x"22" => byteOut <= x"29";
            when x"23" => byteOut <= x"20";
            when x"24" => byteOut <= x"1F";
            when x"25" => byteOut <= x"16";
            when x"26" => byteOut <= x"0D";
            when x"27" => byteOut <= x"04";
            when x"28" => byteOut <= x"73";
            when x"29" => byteOut <= x"7A";
            when x"2A" => byteOut <= x"61";
            when x"2B" => byteOut <= x"68";
            when x"2C" => byteOut <= x"57";
            when x"2D" => byteOut <= x"5E";
            when x"2E" => byteOut <= x"45";
            when x"2F" => byteOut <= x"4C";
            when x"30" => byteOut <= x"AB";
            when x"31" => byteOut <= x"A2";
            when x"32" => byteOut <= x"B9";
            when x"33" => byteOut <= x"B0";
            when x"34" => byteOut <= x"8F";
            when x"35" => byteOut <= x"86";
            when x"36" => byteOut <= x"9D";
            when x"37" => byteOut <= x"94";
            when x"38" => byteOut <= x"E3";
            when x"39" => byteOut <= x"EA";
            when x"3A" => byteOut <= x"F1";
            when x"3B" => byteOut <= x"F8";
            when x"3C" => byteOut <= x"C7";
            when x"3D" => byteOut <= x"CE";
            when x"3E" => byteOut <= x"D5";
            when x"3F" => byteOut <= x"DC";
            when x"40" => byteOut <= x"76";
            when x"41" => byteOut <= x"7F";
            when x"42" => byteOut <= x"64";
            when x"43" => byteOut <= x"6D";
            when x"44" => byteOut <= x"52";
            when x"45" => byteOut <= x"5B";
            when x"46" => byteOut <= x"40";
            when x"47" => byteOut <= x"49";
            when x"48" => byteOut <= x"3E";
            when x"49" => byteOut <= x"37";
            when x"4A" => byteOut <= x"2C";
            when x"4B" => byteOut <= x"25";
            when x"4C" => byteOut <= x"1A";
            when x"4D" => byteOut <= x"13";
            when x"4E" => byteOut <= x"08";
            when x"4F" => byteOut <= x"01";
            when x"50" => byteOut <= x"E6";
            when x"51" => byteOut <= x"EF";
            when x"52" => byteOut <= x"F4";
            when x"53" => byteOut <= x"FD";
            when x"54" => byteOut <= x"C2";
            when x"55" => byteOut <= x"CB";
            when x"56" => byteOut <= x"D0";
            when x"57" => byteOut <= x"D9";
            when x"58" => byteOut <= x"AE";
            when x"59" => byteOut <= x"A7";
            when x"5A" => byteOut <= x"BC";
            when x"5B" => byteOut <= x"B5";
            when x"5C" => byteOut <= x"8A";
            when x"5D" => byteOut <= x"83";
            when x"5E" => byteOut <= x"98";
            when x"5F" => byteOut <= x"91";
            when x"60" => byteOut <= x"4D";
            when x"61" => byteOut <= x"44";
            when x"62" => byteOut <= x"5F";
            when x"63" => byteOut <= x"56";
            when x"64" => byteOut <= x"69";
            when x"65" => byteOut <= x"60";
            when x"66" => byteOut <= x"7B";
            when x"67" => byteOut <= x"72";
            when x"68" => byteOut <= x"05";
            when x"69" => byteOut <= x"0C";
            when x"6A" => byteOut <= x"17";
            when x"6B" => byteOut <= x"1E";
            when x"6C" => byteOut <= x"21";
            when x"6D" => byteOut <= x"28";
            when x"6E" => byteOut <= x"33";
            when x"6F" => byteOut <= x"3A";
            when x"70" => byteOut <= x"DD";
            when x"71" => byteOut <= x"D4";
            when x"72" => byteOut <= x"CF";
            when x"73" => byteOut <= x"C6";
            when x"74" => byteOut <= x"F9";
            when x"75" => byteOut <= x"F0";
            when x"76" => byteOut <= x"EB";
            when x"77" => byteOut <= x"E2";
            when x"78" => byteOut <= x"95";
            when x"79" => byteOut <= x"9C";
            when x"7A" => byteOut <= x"87";
            when x"7B" => byteOut <= x"8E";
            when x"7C" => byteOut <= x"B1";
            when x"7D" => byteOut <= x"B8";
            when x"7E" => byteOut <= x"A3";
            when x"7F" => byteOut <= x"AA";
            when x"80" => byteOut <= x"EC";
            when x"81" => byteOut <= x"E5";
            when x"82" => byteOut <= x"FE";
            when x"83" => byteOut <= x"F7";
            when x"84" => byteOut <= x"C8";
            when x"85" => byteOut <= x"C1";
            when x"86" => byteOut <= x"DA";
            when x"87" => byteOut <= x"D3";
            when x"88" => byteOut <= x"A4";
            when x"89" => byteOut <= x"AD";
            when x"8A" => byteOut <= x"B6";
            when x"8B" => byteOut <= x"BF";
            when x"8C" => byteOut <= x"80";
            when x"8D" => byteOut <= x"89";
            when x"8E" => byteOut <= x"92";
            when x"8F" => byteOut <= x"9B";
            when x"90" => byteOut <= x"7C";
            when x"91" => byteOut <= x"75";
            when x"92" => byteOut <= x"6E";
            when x"93" => byteOut <= x"67";
            when x"94" => byteOut <= x"58";
            when x"95" => byteOut <= x"51";
            when x"96" => byteOut <= x"4A";
            when x"97" => byteOut <= x"43";
            when x"98" => byteOut <= x"34";
            when x"99" => byteOut <= x"3D";
            when x"9A" => byteOut <= x"26";
            when x"9B" => byteOut <= x"2F";
            when x"9C" => byteOut <= x"10";
            when x"9D" => byteOut <= x"19";
            when x"9E" => byteOut <= x"02";
            when x"9F" => byteOut <= x"0B";
            when x"A0" => byteOut <= x"D7";
            when x"A1" => byteOut <= x"DE";
            when x"A2" => byteOut <= x"C5";
            when x"A3" => byteOut <= x"CC";
            when x"A4" => byteOut <= x"F3";
            when x"A5" => byteOut <= x"FA";
            when x"A6" => byteOut <= x"E1";
            when x"A7" => byteOut <= x"E8";
            when x"A8" => byteOut <= x"9F";
            when x"A9" => byteOut <= x"96";
            when x"AA" => byteOut <= x"8D";
            when x"AB" => byteOut <= x"84";
            when x"AC" => byteOut <= x"BB";
            when x"AD" => byteOut <= x"B2";
            when x"AE" => byteOut <= x"A9";
            when x"AF" => byteOut <= x"A0";
            when x"B0" => byteOut <= x"47";
            when x"B1" => byteOut <= x"4E";
            when x"B2" => byteOut <= x"55";
            when x"B3" => byteOut <= x"5C";
            when x"B4" => byteOut <= x"63";
            when x"B5" => byteOut <= x"6A";
            when x"B6" => byteOut <= x"71";
            when x"B7" => byteOut <= x"78";
            when x"B8" => byteOut <= x"0F";
            when x"B9" => byteOut <= x"06";
            when x"BA" => byteOut <= x"1D";
            when x"BB" => byteOut <= x"14";
            when x"BC" => byteOut <= x"2B";
            when x"BD" => byteOut <= x"22";
            when x"BE" => byteOut <= x"39";
            when x"BF" => byteOut <= x"30";
            when x"C0" => byteOut <= x"9A";
            when x"C1" => byteOut <= x"93";
            when x"C2" => byteOut <= x"88";
            when x"C3" => byteOut <= x"81";
            when x"C4" => byteOut <= x"BE";
            when x"C5" => byteOut <= x"B7";
            when x"C6" => byteOut <= x"AC";
            when x"C7" => byteOut <= x"A5";
            when x"C8" => byteOut <= x"D2";
            when x"C9" => byteOut <= x"DB";
            when x"CA" => byteOut <= x"C0";
            when x"CB" => byteOut <= x"C9";
            when x"CC" => byteOut <= x"F6";
            when x"CD" => byteOut <= x"FF";
            when x"CE" => byteOut <= x"E4";
            when x"CF" => byteOut <= x"ED";
            when x"D0" => byteOut <= x"0A";
            when x"D1" => byteOut <= x"03";
            when x"D2" => byteOut <= x"18";
            when x"D3" => byteOut <= x"11";
            when x"D4" => byteOut <= x"2E";
            when x"D5" => byteOut <= x"27";
            when x"D6" => byteOut <= x"3C";
            when x"D7" => byteOut <= x"35";
            when x"D8" => byteOut <= x"42";
            when x"D9" => byteOut <= x"4B";
            when x"DA" => byteOut <= x"50";
            when x"DB" => byteOut <= x"59";
            when x"DC" => byteOut <= x"66";
            when x"DD" => byteOut <= x"6F";
            when x"DE" => byteOut <= x"74";
            when x"DF" => byteOut <= x"7D";
            when x"E0" => byteOut <= x"A1";
            when x"E1" => byteOut <= x"A8";
            when x"E2" => byteOut <= x"B3";
            when x"E3" => byteOut <= x"BA";
            when x"E4" => byteOut <= x"85";
            when x"E5" => byteOut <= x"8C";
            when x"E6" => byteOut <= x"97";
            when x"E7" => byteOut <= x"9E";
            when x"E8" => byteOut <= x"E9";
            when x"E9" => byteOut <= x"E0";
            when x"EA" => byteOut <= x"FB";
            when x"EB" => byteOut <= x"F2";
            when x"EC" => byteOut <= x"CD";
            when x"ED" => byteOut <= x"C4";
            when x"EE" => byteOut <= x"DF";
            when x"EF" => byteOut <= x"D6";
            when x"F0" => byteOut <= x"31";
            when x"F1" => byteOut <= x"38";
            when x"F2" => byteOut <= x"23";
            when x"F3" => byteOut <= x"2A";
            when x"F4" => byteOut <= x"15";
            when x"F5" => byteOut <= x"1C";
            when x"F6" => byteOut <= x"07";
            when x"F7" => byteOut <= x"0E";
            when x"F8" => byteOut <= x"79";
            when x"F9" => byteOut <= x"70";
            when x"FA" => byteOut <= x"6B";
            when x"FB" => byteOut <= x"62";
            when x"FC" => byteOut <= x"5D";
            when x"FD" => byteOut <= x"54";
            when x"FE" => byteOut <= x"4F";
            when x"FF" => byteOut <= x"46";
            when others => byteOut <= x"00";
        end case;
    end process;
end architecture;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity x11 is
    Port ( byteIn : in STD_LOGIC_VECTOR(7 downto 0);
           byteOut : out STD_LOGIC_VECTOR(7 downto 0));
end x11;

architecture Behavioral of x11 is
begin
    process(byteIn)
    begin
        case byteIn is
            when x"00" => byteOut <= x"00";
            when x"01" => byteOut <= x"0B";
            when x"02" => byteOut <= x"16";
            when x"03" => byteOut <= x"1D";
            when x"04" => byteOut <= x"2C";
            when x"05" => byteOut <= x"27";
            when x"06" => byteOut <= x"3A";
            when x"07" => byteOut <= x"31";
            when x"08" => byteOut <= x"58";
            when x"09" => byteOut <= x"53";
            when x"0A" => byteOut <= x"4E";
            when x"0B" => byteOut <= x"45";
            when x"0C" => byteOut <= x"74";
            when x"0D" => byteOut <= x"7F";
            when x"0E" => byteOut <= x"62";
            when x"0F" => byteOut <= x"69";
            when x"10" => byteOut <= x"B0";
            when x"11" => byteOut <= x"BB";
            when x"12" => byteOut <= x"A6";
            when x"13" => byteOut <= x"AD";
            when x"14" => byteOut <= x"9C";
            when x"15" => byteOut <= x"97";
            when x"16" => byteOut <= x"8A";
            when x"17" => byteOut <= x"81";
            when x"18" => byteOut <= x"E8";
            when x"19" => byteOut <= x"E3";
            when x"1A" => byteOut <= x"FE";
            when x"1B" => byteOut <= x"F5";
            when x"1C" => byteOut <= x"C4";
            when x"1D" => byteOut <= x"CF";
            when x"1E" => byteOut <= x"D2";
            when x"1F" => byteOut <= x"D9";
            when x"20" => byteOut <= x"7B";
            when x"21" => byteOut <= x"70";
            when x"22" => byteOut <= x"6D";
            when x"23" => byteOut <= x"66";
            when x"24" => byteOut <= x"57";
            when x"25" => byteOut <= x"5C";
            when x"26" => byteOut <= x"41";
            when x"27" => byteOut <= x"4A";
            when x"28" => byteOut <= x"23";
            when x"29" => byteOut <= x"28";
            when x"2A" => byteOut <= x"35";
            when x"2B" => byteOut <= x"3E";
            when x"2C" => byteOut <= x"0F";
            when x"2D" => byteOut <= x"04";
            when x"2E" => byteOut <= x"19";
            when x"2F" => byteOut <= x"12";
            when x"30" => byteOut <= x"CB";
            when x"31" => byteOut <= x"C0";
            when x"32" => byteOut <= x"DD";
            when x"33" => byteOut <= x"D6";
            when x"34" => byteOut <= x"E7";
            when x"35" => byteOut <= x"EC";
            when x"36" => byteOut <= x"F1";
            when x"37" => byteOut <= x"FA";
            when x"38" => byteOut <= x"93";
            when x"39" => byteOut <= x"98";
            when x"3A" => byteOut <= x"85";
            when x"3B" => byteOut <= x"8E";
            when x"3C" => byteOut <= x"BF";
            when x"3D" => byteOut <= x"B4";
            when x"3E" => byteOut <= x"A9";
            when x"3F" => byteOut <= x"A2";
            when x"40" => byteOut <= x"F6";
            when x"41" => byteOut <= x"FD";
            when x"42" => byteOut <= x"E0";
            when x"43" => byteOut <= x"EB";
            when x"44" => byteOut <= x"DA";
            when x"45" => byteOut <= x"D1";
            when x"46" => byteOut <= x"CC";
            when x"47" => byteOut <= x"C7";
            when x"48" => byteOut <= x"AE";
            when x"49" => byteOut <= x"A5";
            when x"4A" => byteOut <= x"B8";
            when x"4B" => byteOut <= x"B3";
            when x"4C" => byteOut <= x"82";
            when x"4D" => byteOut <= x"89";
            when x"4E" => byteOut <= x"94";
            when x"4F" => byteOut <= x"9F";
            when x"50" => byteOut <= x"46";
            when x"51" => byteOut <= x"4D";
            when x"52" => byteOut <= x"50";
            when x"53" => byteOut <= x"5B";
            when x"54" => byteOut <= x"6A";
            when x"55" => byteOut <= x"61";
            when x"56" => byteOut <= x"7C";
            when x"57" => byteOut <= x"77";
            when x"58" => byteOut <= x"1E";
            when x"59" => byteOut <= x"15";
            when x"5A" => byteOut <= x"08";
            when x"5B" => byteOut <= x"03";
            when x"5C" => byteOut <= x"32";
            when x"5D" => byteOut <= x"39";
            when x"5E" => byteOut <= x"24";
            when x"5F" => byteOut <= x"2F";
            when x"60" => byteOut <= x"8D";
            when x"61" => byteOut <= x"86";
            when x"62" => byteOut <= x"9B";
            when x"63" => byteOut <= x"90";
            when x"64" => byteOut <= x"A1";
            when x"65" => byteOut <= x"AA";
            when x"66" => byteOut <= x"B7";
            when x"67" => byteOut <= x"BC";
            when x"68" => byteOut <= x"D5";
            when x"69" => byteOut <= x"DE";
            when x"6A" => byteOut <= x"C3";
            when x"6B" => byteOut <= x"C8";
            when x"6C" => byteOut <= x"F9";
            when x"6D" => byteOut <= x"F2";
            when x"6E" => byteOut <= x"EF";
            when x"6F" => byteOut <= x"E4";
            when x"70" => byteOut <= x"3D";
            when x"71" => byteOut <= x"36";
            when x"72" => byteOut <= x"2B";
            when x"73" => byteOut <= x"20";
            when x"74" => byteOut <= x"11";
            when x"75" => byteOut <= x"1A";
            when x"76" => byteOut <= x"07";
            when x"77" => byteOut <= x"0C";
            when x"78" => byteOut <= x"65";
            when x"79" => byteOut <= x"6E";
            when x"7A" => byteOut <= x"73";
            when x"7B" => byteOut <= x"78";
            when x"7C" => byteOut <= x"49";
            when x"7D" => byteOut <= x"42";
            when x"7E" => byteOut <= x"5F";
            when x"7F" => byteOut <= x"54";
            when x"80" => byteOut <= x"F7";
            when x"81" => byteOut <= x"FC";
            when x"82" => byteOut <= x"E1";
            when x"83" => byteOut <= x"EA";
            when x"84" => byteOut <= x"DB";
            when x"85" => byteOut <= x"D0";
            when x"86" => byteOut <= x"CD";
            when x"87" => byteOut <= x"C6";
            when x"88" => byteOut <= x"AF";
            when x"89" => byteOut <= x"A4";
            when x"8A" => byteOut <= x"B9";
            when x"8B" => byteOut <= x"B2";
            when x"8C" => byteOut <= x"83";
            when x"8D" => byteOut <= x"88";
            when x"8E" => byteOut <= x"95";
            when x"8F" => byteOut <= x"9E";
            when x"90" => byteOut <= x"47";
            when x"91" => byteOut <= x"4C";
            when x"92" => byteOut <= x"51";
            when x"93" => byteOut <= x"5A";
            when x"94" => byteOut <= x"6B";
            when x"95" => byteOut <= x"60";
            when x"96" => byteOut <= x"7D";
            when x"97" => byteOut <= x"76";
            when x"98" => byteOut <= x"1F";
            when x"99" => byteOut <= x"14";
            when x"9A" => byteOut <= x"09";
            when x"9B" => byteOut <= x"02";
            when x"9C" => byteOut <= x"33";
            when x"9D" => byteOut <= x"38";
            when x"9E" => byteOut <= x"25";
            when x"9F" => byteOut <= x"2E";
            when x"A0" => byteOut <= x"8C";
            when x"A1" => byteOut <= x"87";
            when x"A2" => byteOut <= x"9A";
            when x"A3" => byteOut <= x"91";
            when x"A4" => byteOut <= x"A0";
            when x"A5" => byteOut <= x"AB";
            when x"A6" => byteOut <= x"B6";
            when x"A7" => byteOut <= x"BD";
            when x"A8" => byteOut <= x"D4";
            when x"A9" => byteOut <= x"DF";
            when x"AA" => byteOut <= x"C2";
            when x"AB" => byteOut <= x"C9";
            when x"AC" => byteOut <= x"F8";
            when x"AD" => byteOut <= x"F3";
            when x"AE" => byteOut <= x"EE";
            when x"AF" => byteOut <= x"E5";
            when x"B0" => byteOut <= x"3C";
            when x"B1" => byteOut <= x"37";
            when x"B2" => byteOut <= x"2A";
            when x"B3" => byteOut <= x"21";
            when x"B4" => byteOut <= x"10";
            when x"B5" => byteOut <= x"1B";
            when x"B6" => byteOut <= x"06";
            when x"B7" => byteOut <= x"0D";
            when x"B8" => byteOut <= x"64";
            when x"B9" => byteOut <= x"6F";
            when x"BA" => byteOut <= x"72";
            when x"BB" => byteOut <= x"79";
            when x"BC" => byteOut <= x"48";
            when x"BD" => byteOut <= x"43";
            when x"BE" => byteOut <= x"5E";
            when x"BF" => byteOut <= x"55";
            when x"C0" => byteOut <= x"01";
            when x"C1" => byteOut <= x"0A";
            when x"C2" => byteOut <= x"17";
            when x"C3" => byteOut <= x"1C";
            when x"C4" => byteOut <= x"2D";
            when x"C5" => byteOut <= x"26";
            when x"C6" => byteOut <= x"3B";
            when x"C7" => byteOut <= x"30";
            when x"C8" => byteOut <= x"59";
            when x"C9" => byteOut <= x"52";
            when x"CA" => byteOut <= x"4F";
            when x"CB" => byteOut <= x"44";
            when x"CC" => byteOut <= x"75";
            when x"CD" => byteOut <= x"7E";
            when x"CE" => byteOut <= x"63";
            when x"CF" => byteOut <= x"68";
            when x"D0" => byteOut <= x"B1";
            when x"D1" => byteOut <= x"BA";
            when x"D2" => byteOut <= x"A7";
            when x"D3" => byteOut <= x"AC";
            when x"D4" => byteOut <= x"9D";
            when x"D5" => byteOut <= x"96";
            when x"D6" => byteOut <= x"8B";
            when x"D7" => byteOut <= x"80";
            when x"D8" => byteOut <= x"E9";
            when x"D9" => byteOut <= x"E2";
            when x"DA" => byteOut <= x"FF";
            when x"DB" => byteOut <= x"F4";
            when x"DC" => byteOut <= x"C5";
            when x"DD" => byteOut <= x"CE";
            when x"DE" => byteOut <= x"D3";
            when x"DF" => byteOut <= x"D8";
            when x"E0" => byteOut <= x"7A";
            when x"E1" => byteOut <= x"71";
            when x"E2" => byteOut <= x"6C";
            when x"E3" => byteOut <= x"67";
            when x"E4" => byteOut <= x"56";
            when x"E5" => byteOut <= x"5D";
            when x"E6" => byteOut <= x"40";
            when x"E7" => byteOut <= x"4B";
            when x"E8" => byteOut <= x"22";
            when x"E9" => byteOut <= x"29";
            when x"EA" => byteOut <= x"34";
            when x"EB" => byteOut <= x"3F";
            when x"EC" => byteOut <= x"0E";
            when x"ED" => byteOut <= x"05";
            when x"EE" => byteOut <= x"18";
            when x"EF" => byteOut <= x"13";
            when x"F0" => byteOut <= x"CA";
            when x"F1" => byteOut <= x"C1";
            when x"F2" => byteOut <= x"DC";
            when x"F3" => byteOut <= x"D7";
            when x"F4" => byteOut <= x"E6";
            when x"F5" => byteOut <= x"ED";
            when x"F6" => byteOut <= x"F0";
            when x"F7" => byteOut <= x"FB";
            when x"F8" => byteOut <= x"92";
            when x"F9" => byteOut <= x"99";
            when x"FA" => byteOut <= x"84";
            when x"FB" => byteOut <= x"8F";
            when x"FC" => byteOut <= x"BE";
            when x"FD" => byteOut <= x"B5";
            when x"FE" => byteOut <= x"A8";
            when x"FF" => byteOut <= x"A3";
            when others => byteOut <= x"00";
        end case;
    end process;
end architecture;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity x13 is
    Port ( byteIn : in STD_LOGIC_VECTOR(7 downto 0);
           byteOut : out STD_LOGIC_VECTOR(7 downto 0));
end x13;

architecture Behavioral of x13 is
begin
    process(byteIn)
    begin
        case byteIn is
            when x"00" => byteOut <= x"00";
            when x"01" => byteOut <= x"0D";
            when x"02" => byteOut <= x"1A";
            when x"03" => byteOut <= x"17";
            when x"04" => byteOut <= x"34";
            when x"05" => byteOut <= x"39";
            when x"06" => byteOut <= x"2E";
            when x"07" => byteOut <= x"23";
            when x"08" => byteOut <= x"68";
            when x"09" => byteOut <= x"65";
            when x"0A" => byteOut <= x"72";
            when x"0B" => byteOut <= x"7F";
            when x"0C" => byteOut <= x"5C";
            when x"0D" => byteOut <= x"51";
            when x"0E" => byteOut <= x"46";
            when x"0F" => byteOut <= x"4B";
            when x"10" => byteOut <= x"D0";
            when x"11" => byteOut <= x"DD";
            when x"12" => byteOut <= x"CA";
            when x"13" => byteOut <= x"C7";
            when x"14" => byteOut <= x"E4";
            when x"15" => byteOut <= x"E9";
            when x"16" => byteOut <= x"FE";
            when x"17" => byteOut <= x"F3";
            when x"18" => byteOut <= x"B8";
            when x"19" => byteOut <= x"B5";
            when x"1A" => byteOut <= x"A2";
            when x"1B" => byteOut <= x"AF";
            when x"1C" => byteOut <= x"8C";
            when x"1D" => byteOut <= x"81";
            when x"1E" => byteOut <= x"96";
            when x"1F" => byteOut <= x"9B";
            when x"20" => byteOut <= x"BB";
            when x"21" => byteOut <= x"B6";
            when x"22" => byteOut <= x"A1";
            when x"23" => byteOut <= x"AC";
            when x"24" => byteOut <= x"8F";
            when x"25" => byteOut <= x"82";
            when x"26" => byteOut <= x"95";
            when x"27" => byteOut <= x"98";
            when x"28" => byteOut <= x"D3";
            when x"29" => byteOut <= x"DE";
            when x"2A" => byteOut <= x"C9";
            when x"2B" => byteOut <= x"C4";
            when x"2C" => byteOut <= x"E7";
            when x"2D" => byteOut <= x"EA";
            when x"2E" => byteOut <= x"FD";
            when x"2F" => byteOut <= x"F0";
            when x"30" => byteOut <= x"6B";
            when x"31" => byteOut <= x"66";
            when x"32" => byteOut <= x"71";
            when x"33" => byteOut <= x"7C";
            when x"34" => byteOut <= x"5F";
            when x"35" => byteOut <= x"52";
            when x"36" => byteOut <= x"45";
            when x"37" => byteOut <= x"48";
            when x"38" => byteOut <= x"03";
            when x"39" => byteOut <= x"0E";
            when x"3A" => byteOut <= x"19";
            when x"3B" => byteOut <= x"14";
            when x"3C" => byteOut <= x"37";
            when x"3D" => byteOut <= x"3A";
            when x"3E" => byteOut <= x"2D";
            when x"3F" => byteOut <= x"20";
            when x"40" => byteOut <= x"6D";
            when x"41" => byteOut <= x"60";
            when x"42" => byteOut <= x"77";
            when x"43" => byteOut <= x"7A";
            when x"44" => byteOut <= x"59";
            when x"45" => byteOut <= x"54";
            when x"46" => byteOut <= x"43";
            when x"47" => byteOut <= x"4E";
            when x"48" => byteOut <= x"05";
            when x"49" => byteOut <= x"08";
            when x"4A" => byteOut <= x"1F";
            when x"4B" => byteOut <= x"12";
            when x"4C" => byteOut <= x"31";
            when x"4D" => byteOut <= x"3C";
            when x"4E" => byteOut <= x"2B";
            when x"4F" => byteOut <= x"26";
            when x"50" => byteOut <= x"BD";
            when x"51" => byteOut <= x"B0";
            when x"52" => byteOut <= x"A7";
            when x"53" => byteOut <= x"AA";
            when x"54" => byteOut <= x"89";
            when x"55" => byteOut <= x"84";
            when x"56" => byteOut <= x"93";
            when x"57" => byteOut <= x"9E";
            when x"58" => byteOut <= x"D5";
            when x"59" => byteOut <= x"D8";
            when x"5A" => byteOut <= x"CF";
            when x"5B" => byteOut <= x"C2";
            when x"5C" => byteOut <= x"E1";
            when x"5D" => byteOut <= x"EC";
            when x"5E" => byteOut <= x"FB";
            when x"5F" => byteOut <= x"F6";
            when x"60" => byteOut <= x"D6";
            when x"61" => byteOut <= x"DB";
            when x"62" => byteOut <= x"CC";
            when x"63" => byteOut <= x"C1";
            when x"64" => byteOut <= x"E2";
            when x"65" => byteOut <= x"EF";
            when x"66" => byteOut <= x"F8";
            when x"67" => byteOut <= x"F5";
            when x"68" => byteOut <= x"BE";
            when x"69" => byteOut <= x"B3";
            when x"6A" => byteOut <= x"A4";
            when x"6B" => byteOut <= x"A9";
            when x"6C" => byteOut <= x"8A";
            when x"6D" => byteOut <= x"87";
            when x"6E" => byteOut <= x"90";
            when x"6F" => byteOut <= x"9D";
            when x"70" => byteOut <= x"06";
            when x"71" => byteOut <= x"0B";
            when x"72" => byteOut <= x"1C";
            when x"73" => byteOut <= x"11";
            when x"74" => byteOut <= x"32";
            when x"75" => byteOut <= x"3F";
            when x"76" => byteOut <= x"28";
            when x"77" => byteOut <= x"25";
            when x"78" => byteOut <= x"6E";
            when x"79" => byteOut <= x"63";
            when x"7A" => byteOut <= x"74";
            when x"7B" => byteOut <= x"79";
            when x"7C" => byteOut <= x"5A";
            when x"7D" => byteOut <= x"57";
            when x"7E" => byteOut <= x"40";
            when x"7F" => byteOut <= x"4D";
            when x"80" => byteOut <= x"DA";
            when x"81" => byteOut <= x"D7";
            when x"82" => byteOut <= x"C0";
            when x"83" => byteOut <= x"CD";
            when x"84" => byteOut <= x"EE";
            when x"85" => byteOut <= x"E3";
            when x"86" => byteOut <= x"F4";
            when x"87" => byteOut <= x"F9";
            when x"88" => byteOut <= x"B2";
            when x"89" => byteOut <= x"BF";
            when x"8A" => byteOut <= x"A8";
            when x"8B" => byteOut <= x"A5";
            when x"8C" => byteOut <= x"86";
            when x"8D" => byteOut <= x"8B";
            when x"8E" => byteOut <= x"9C";
            when x"8F" => byteOut <= x"91";
            when x"90" => byteOut <= x"0A";
            when x"91" => byteOut <= x"07";
            when x"92" => byteOut <= x"10";
            when x"93" => byteOut <= x"1D";
            when x"94" => byteOut <= x"3E";
            when x"95" => byteOut <= x"33";
            when x"96" => byteOut <= x"24";
            when x"97" => byteOut <= x"29";
            when x"98" => byteOut <= x"62";
            when x"99" => byteOut <= x"6F";
            when x"9A" => byteOut <= x"78";
            when x"9B" => byteOut <= x"75";
            when x"9C" => byteOut <= x"56";
            when x"9D" => byteOut <= x"5B";
            when x"9E" => byteOut <= x"4C";
            when x"9F" => byteOut <= x"41";
            when x"A0" => byteOut <= x"61";
            when x"A1" => byteOut <= x"6C";
            when x"A2" => byteOut <= x"7B";
            when x"A3" => byteOut <= x"76";
            when x"A4" => byteOut <= x"55";
            when x"A5" => byteOut <= x"58";
            when x"A6" => byteOut <= x"4F";
            when x"A7" => byteOut <= x"42";
            when x"A8" => byteOut <= x"09";
            when x"A9" => byteOut <= x"04";
            when x"AA" => byteOut <= x"13";
            when x"AB" => byteOut <= x"1E";
            when x"AC" => byteOut <= x"3D";
            when x"AD" => byteOut <= x"30";
            when x"AE" => byteOut <= x"27";
            when x"AF" => byteOut <= x"2A";
            when x"B0" => byteOut <= x"B1";
            when x"B1" => byteOut <= x"BC";
            when x"B2" => byteOut <= x"AB";
            when x"B3" => byteOut <= x"A6";
            when x"B4" => byteOut <= x"85";
            when x"B5" => byteOut <= x"88";
            when x"B6" => byteOut <= x"9F";
            when x"B7" => byteOut <= x"92";
            when x"B8" => byteOut <= x"D9";
            when x"B9" => byteOut <= x"D4";
            when x"BA" => byteOut <= x"C3";
            when x"BB" => byteOut <= x"CE";
            when x"BC" => byteOut <= x"ED";
            when x"BD" => byteOut <= x"E0";
            when x"BE" => byteOut <= x"F7";
            when x"BF" => byteOut <= x"FA";
            when x"C0" => byteOut <= x"B7";
            when x"C1" => byteOut <= x"BA";
            when x"C2" => byteOut <= x"AD";
            when x"C3" => byteOut <= x"A0";
            when x"C4" => byteOut <= x"83";
            when x"C5" => byteOut <= x"8E";
            when x"C6" => byteOut <= x"99";
            when x"C7" => byteOut <= x"94";
            when x"C8" => byteOut <= x"DF";
            when x"C9" => byteOut <= x"D2";
            when x"CA" => byteOut <= x"C5";
            when x"CB" => byteOut <= x"C8";
            when x"CC" => byteOut <= x"EB";
            when x"CD" => byteOut <= x"E6";
            when x"CE" => byteOut <= x"F1";
            when x"CF" => byteOut <= x"FC";
            when x"D0" => byteOut <= x"67";
            when x"D1" => byteOut <= x"6A";
            when x"D2" => byteOut <= x"7D";
            when x"D3" => byteOut <= x"70";
            when x"D4" => byteOut <= x"53";
            when x"D5" => byteOut <= x"5E";
            when x"D6" => byteOut <= x"49";
            when x"D7" => byteOut <= x"44";
            when x"D8" => byteOut <= x"0F";
            when x"D9" => byteOut <= x"02";
            when x"DA" => byteOut <= x"15";
            when x"DB" => byteOut <= x"18";
            when x"DC" => byteOut <= x"3B";
            when x"DD" => byteOut <= x"36";
            when x"DE" => byteOut <= x"21";
            when x"DF" => byteOut <= x"2C";
            when x"E0" => byteOut <= x"0C";
            when x"E1" => byteOut <= x"01";
            when x"E2" => byteOut <= x"16";
            when x"E3" => byteOut <= x"1B";
            when x"E4" => byteOut <= x"38";
            when x"E5" => byteOut <= x"35";
            when x"E6" => byteOut <= x"22";
            when x"E7" => byteOut <= x"2F";
            when x"E8" => byteOut <= x"64";
            when x"E9" => byteOut <= x"69";
            when x"EA" => byteOut <= x"7E";
            when x"EB" => byteOut <= x"73";
            when x"EC" => byteOut <= x"50";
            when x"ED" => byteOut <= x"5D";
            when x"EE" => byteOut <= x"4A";
            when x"EF" => byteOut <= x"47";
            when x"F0" => byteOut <= x"DC";
            when x"F1" => byteOut <= x"D1";
            when x"F2" => byteOut <= x"C6";
            when x"F3" => byteOut <= x"CB";
            when x"F4" => byteOut <= x"E8";
            when x"F5" => byteOut <= x"E5";
            when x"F6" => byteOut <= x"F2";
            when x"F7" => byteOut <= x"FF";
            when x"F8" => byteOut <= x"B4";
            when x"F9" => byteOut <= x"B9";
            when x"FA" => byteOut <= x"AE";
            when x"FB" => byteOut <= x"A3";
            when x"FC" => byteOut <= x"80";
            when x"FD" => byteOut <= x"8D";
            when x"FE" => byteOut <= x"9A";
            when x"FF" => byteOut <= x"97";
            when others => byteOut <= x"00";
        end case;
    end process;
end architecture;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity x14 is
    Port ( byteIn : in STD_LOGIC_VECTOR(7 downto 0);
           byteOut : out STD_LOGIC_VECTOR(7 downto 0));
end x14;

architecture Behavioral of x14 is
begin
    process(byteIn)
    begin
        case byteIn is
            when x"00" => byteOut <= x"00";
            when x"01" => byteOut <= x"0E";
            when x"02" => byteOut <= x"1C";
            when x"03" => byteOut <= x"12";
            when x"04" => byteOut <= x"38";
            when x"05" => byteOut <= x"36";
            when x"06" => byteOut <= x"24";
            when x"07" => byteOut <= x"2A";
            when x"08" => byteOut <= x"70";
            when x"09" => byteOut <= x"7E";
            when x"0A" => byteOut <= x"6C";
            when x"0B" => byteOut <= x"62";
            when x"0C" => byteOut <= x"48";
            when x"0D" => byteOut <= x"46";
            when x"0E" => byteOut <= x"54";
            when x"0F" => byteOut <= x"5A";
            when x"10" => byteOut <= x"E0";
            when x"11" => byteOut <= x"EE";
            when x"12" => byteOut <= x"FC";
            when x"13" => byteOut <= x"F2";
            when x"14" => byteOut <= x"D8";
            when x"15" => byteOut <= x"D6";
            when x"16" => byteOut <= x"C4";
            when x"17" => byteOut <= x"CA";
            when x"18" => byteOut <= x"90";
            when x"19" => byteOut <= x"9E";
            when x"1A" => byteOut <= x"8C";
            when x"1B" => byteOut <= x"82";
            when x"1C" => byteOut <= x"A8";
            when x"1D" => byteOut <= x"A6";
            when x"1E" => byteOut <= x"B4";
            when x"1F" => byteOut <= x"BA";
            when x"20" => byteOut <= x"DB";
            when x"21" => byteOut <= x"D5";
            when x"22" => byteOut <= x"C7";
            when x"23" => byteOut <= x"C9";
            when x"24" => byteOut <= x"E3";
            when x"25" => byteOut <= x"ED";
            when x"26" => byteOut <= x"FF";
            when x"27" => byteOut <= x"F1";
            when x"28" => byteOut <= x"AB";
            when x"29" => byteOut <= x"A5";
            when x"2A" => byteOut <= x"B7";
            when x"2B" => byteOut <= x"B9";
            when x"2C" => byteOut <= x"93";
            when x"2D" => byteOut <= x"9D";
            when x"2E" => byteOut <= x"8F";
            when x"2F" => byteOut <= x"81";
            when x"30" => byteOut <= x"3B";
            when x"31" => byteOut <= x"35";
            when x"32" => byteOut <= x"27";
            when x"33" => byteOut <= x"29";
            when x"34" => byteOut <= x"03";
            when x"35" => byteOut <= x"0D";
            when x"36" => byteOut <= x"1F";
            when x"37" => byteOut <= x"11";
            when x"38" => byteOut <= x"4B";
            when x"39" => byteOut <= x"45";
            when x"3A" => byteOut <= x"57";
            when x"3B" => byteOut <= x"59";
            when x"3C" => byteOut <= x"73";
            when x"3D" => byteOut <= x"7D";
            when x"3E" => byteOut <= x"6F";
            when x"3F" => byteOut <= x"61";
            when x"40" => byteOut <= x"AD";
            when x"41" => byteOut <= x"A3";
            when x"42" => byteOut <= x"B1";
            when x"43" => byteOut <= x"BF";
            when x"44" => byteOut <= x"95";
            when x"45" => byteOut <= x"9B";
            when x"46" => byteOut <= x"89";
            when x"47" => byteOut <= x"87";
            when x"48" => byteOut <= x"DD";
            when x"49" => byteOut <= x"D3";
            when x"4A" => byteOut <= x"C1";
            when x"4B" => byteOut <= x"CF";
            when x"4C" => byteOut <= x"E5";
            when x"4D" => byteOut <= x"EB";
            when x"4E" => byteOut <= x"F9";
            when x"4F" => byteOut <= x"F7";
            when x"50" => byteOut <= x"4D";
            when x"51" => byteOut <= x"43";
            when x"52" => byteOut <= x"51";
            when x"53" => byteOut <= x"5F";
            when x"54" => byteOut <= x"75";
            when x"55" => byteOut <= x"7B";
            when x"56" => byteOut <= x"69";
            when x"57" => byteOut <= x"67";
            when x"58" => byteOut <= x"3D";
            when x"59" => byteOut <= x"33";
            when x"5A" => byteOut <= x"21";
            when x"5B" => byteOut <= x"2F";
            when x"5C" => byteOut <= x"05";
            when x"5D" => byteOut <= x"0B";
            when x"5E" => byteOut <= x"19";
            when x"5F" => byteOut <= x"17";
            when x"60" => byteOut <= x"76";
            when x"61" => byteOut <= x"78";
            when x"62" => byteOut <= x"6A";
            when x"63" => byteOut <= x"64";
            when x"64" => byteOut <= x"4E";
            when x"65" => byteOut <= x"40";
            when x"66" => byteOut <= x"52";
            when x"67" => byteOut <= x"5C";
            when x"68" => byteOut <= x"06";
            when x"69" => byteOut <= x"08";
            when x"6A" => byteOut <= x"1A";
            when x"6B" => byteOut <= x"14";
            when x"6C" => byteOut <= x"3E";
            when x"6D" => byteOut <= x"30";
            when x"6E" => byteOut <= x"22";
            when x"6F" => byteOut <= x"2C";
            when x"70" => byteOut <= x"96";
            when x"71" => byteOut <= x"98";
            when x"72" => byteOut <= x"8A";
            when x"73" => byteOut <= x"84";
            when x"74" => byteOut <= x"AE";
            when x"75" => byteOut <= x"A0";
            when x"76" => byteOut <= x"B2";
            when x"77" => byteOut <= x"BC";
            when x"78" => byteOut <= x"E6";
            when x"79" => byteOut <= x"E8";
            when x"7A" => byteOut <= x"FA";
            when x"7B" => byteOut <= x"F4";
            when x"7C" => byteOut <= x"DE";
            when x"7D" => byteOut <= x"D0";
            when x"7E" => byteOut <= x"C2";
            when x"7F" => byteOut <= x"CC";
            when x"80" => byteOut <= x"41";
            when x"81" => byteOut <= x"4F";
            when x"82" => byteOut <= x"5D";
            when x"83" => byteOut <= x"53";
            when x"84" => byteOut <= x"79";
            when x"85" => byteOut <= x"77";
            when x"86" => byteOut <= x"65";
            when x"87" => byteOut <= x"6B";
            when x"88" => byteOut <= x"31";
            when x"89" => byteOut <= x"3F";
            when x"8A" => byteOut <= x"2D";
            when x"8B" => byteOut <= x"23";
            when x"8C" => byteOut <= x"09";
            when x"8D" => byteOut <= x"07";
            when x"8E" => byteOut <= x"15";
            when x"8F" => byteOut <= x"1B";
            when x"90" => byteOut <= x"A1";
            when x"91" => byteOut <= x"AF";
            when x"92" => byteOut <= x"BD";
            when x"93" => byteOut <= x"B3";
            when x"94" => byteOut <= x"99";
            when x"95" => byteOut <= x"97";
            when x"96" => byteOut <= x"85";
            when x"97" => byteOut <= x"8B";
            when x"98" => byteOut <= x"D1";
            when x"99" => byteOut <= x"DF";
            when x"9A" => byteOut <= x"CD";
            when x"9B" => byteOut <= x"C3";
            when x"9C" => byteOut <= x"E9";
            when x"9D" => byteOut <= x"E7";
            when x"9E" => byteOut <= x"F5";
            when x"9F" => byteOut <= x"FB";
            when x"A0" => byteOut <= x"9A";
            when x"A1" => byteOut <= x"94";
            when x"A2" => byteOut <= x"86";
            when x"A3" => byteOut <= x"88";
            when x"A4" => byteOut <= x"A2";
            when x"A5" => byteOut <= x"AC";
            when x"A6" => byteOut <= x"BE";
            when x"A7" => byteOut <= x"B0";
            when x"A8" => byteOut <= x"EA";
            when x"A9" => byteOut <= x"E4";
            when x"AA" => byteOut <= x"F6";
            when x"AB" => byteOut <= x"F8";
            when x"AC" => byteOut <= x"D2";
            when x"AD" => byteOut <= x"DC";
            when x"AE" => byteOut <= x"CE";
            when x"AF" => byteOut <= x"C0";
            when x"B0" => byteOut <= x"7A";
            when x"B1" => byteOut <= x"74";
            when x"B2" => byteOut <= x"66";
            when x"B3" => byteOut <= x"68";
            when x"B4" => byteOut <= x"42";
            when x"B5" => byteOut <= x"4C";
            when x"B6" => byteOut <= x"5E";
            when x"B7" => byteOut <= x"50";
            when x"B8" => byteOut <= x"0A";
            when x"B9" => byteOut <= x"04";
            when x"BA" => byteOut <= x"16";
            when x"BB" => byteOut <= x"18";
            when x"BC" => byteOut <= x"32";
            when x"BD" => byteOut <= x"3C";
            when x"BE" => byteOut <= x"2E";
            when x"BF" => byteOut <= x"20";
            when x"C0" => byteOut <= x"EC";
            when x"C1" => byteOut <= x"E2";
            when x"C2" => byteOut <= x"F0";
            when x"C3" => byteOut <= x"FE";
            when x"C4" => byteOut <= x"D4";
            when x"C5" => byteOut <= x"DA";
            when x"C6" => byteOut <= x"C8";
            when x"C7" => byteOut <= x"C6";
            when x"C8" => byteOut <= x"9C";
            when x"C9" => byteOut <= x"92";
            when x"CA" => byteOut <= x"80";
            when x"CB" => byteOut <= x"8E";
            when x"CC" => byteOut <= x"A4";
            when x"CD" => byteOut <= x"AA";
            when x"CE" => byteOut <= x"B8";
            when x"CF" => byteOut <= x"B6";
            when x"D0" => byteOut <= x"0C";
            when x"D1" => byteOut <= x"02";
            when x"D2" => byteOut <= x"10";
            when x"D3" => byteOut <= x"1E";
            when x"D4" => byteOut <= x"34";
            when x"D5" => byteOut <= x"3A";
            when x"D6" => byteOut <= x"28";
            when x"D7" => byteOut <= x"26";
            when x"D8" => byteOut <= x"7C";
            when x"D9" => byteOut <= x"72";
            when x"DA" => byteOut <= x"60";
            when x"DB" => byteOut <= x"6E";
            when x"DC" => byteOut <= x"44";
            when x"DD" => byteOut <= x"4A";
            when x"DE" => byteOut <= x"58";
            when x"DF" => byteOut <= x"56";
            when x"E0" => byteOut <= x"37";
            when x"E1" => byteOut <= x"39";
            when x"E2" => byteOut <= x"2B";
            when x"E3" => byteOut <= x"25";
            when x"E4" => byteOut <= x"0F";
            when x"E5" => byteOut <= x"01";
            when x"E6" => byteOut <= x"13";
            when x"E7" => byteOut <= x"1D";
            when x"E8" => byteOut <= x"47";
            when x"E9" => byteOut <= x"49";
            when x"EA" => byteOut <= x"5B";
            when x"EB" => byteOut <= x"55";
            when x"EC" => byteOut <= x"7F";
            when x"ED" => byteOut <= x"71";
            when x"EE" => byteOut <= x"63";
            when x"EF" => byteOut <= x"6D";
            when x"F0" => byteOut <= x"D7";
            when x"F1" => byteOut <= x"D9";
            when x"F2" => byteOut <= x"CB";
            when x"F3" => byteOut <= x"C5";
            when x"F4" => byteOut <= x"EF";
            when x"F5" => byteOut <= x"E1";
            when x"F6" => byteOut <= x"F3";
            when x"F7" => byteOut <= x"FD";
            when x"F8" => byteOut <= x"A7";
            when x"F9" => byteOut <= x"A9";
            when x"FA" => byteOut <= x"BB";
            when x"FB" => byteOut <= x"B5";
            when x"FC" => byteOut <= x"9F";
            when x"FD" => byteOut <= x"91";
            when x"FE" => byteOut <= x"83";
            when x"FF" => byteOut <= x"8D";
            when others => byteOut <= x"00";
        end case;
    end process;
end architecture;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity invMixColumn is
    Port ( wordIn : in STD_LOGIC_VECTOR (31 downto 0);
           wordOut : out STD_LOGIC_VECTOR (31 downto 0));
end invMixColumn;

architecture Behavioral of invMixColumn is
    signal t0_x1, t0_x9, t0_x11, t0_x13, t0_x14 : STD_LOGIC_VECTOR(7 downto 0);
    signal t1_x1, t1_x9, t1_x11, t1_x13, t1_x14 : STD_LOGIC_VECTOR(7 downto 0);
    signal t2_x1, t2_x9, t2_x11, t2_x13, t2_x14 : STD_LOGIC_VECTOR(7 downto 0);
    signal t3_x1, t3_x9, t3_x11, t3_x13, t3_x14 : STD_LOGIC_VECTOR(7 downto 0);
    
    component x9
        Port ( byteIn : in STD_LOGIC_VECTOR(7 downto 0);
               byteOut : out STD_LOGIC_VECTOR(7 downto 0));
    end component;
    
    component x11
        Port ( byteIn : in STD_LOGIC_VECTOR(7 downto 0);
               byteOut : out STD_LOGIC_VECTOR(7 downto 0));
    end component;
        
    component x13
        Port ( byteIn : in STD_LOGIC_VECTOR(7 downto 0);
               byteOut : out STD_LOGIC_VECTOR(7 downto 0));
    end component;
            
    component x14
        Port ( byteIn : in STD_LOGIC_VECTOR(7 downto 0);
               byteOut : out STD_LOGIC_VECTOR(7 downto 0));
    end component;
begin
    t0_x1 <= wordIn(31 downto 24);
    t1_x1 <= wordIn(23 downto 16);
    t2_x1 <= wordIn(15 downto 8);
    t3_x1 <= wordIn(7 downto 0);
    
    t0x9: x9 port map(byteIn => t0_x1, byteOut => t0_x9);
    t1x9: x9 port map(byteIn => t1_x1, byteOut => t1_x9);
    t2x9: x9 port map(byteIn => t2_x1, byteOut => t2_x9);
    t3x9: x9 port map(byteIn => t3_x1, byteOut => t3_x9);

    t0x11: x11 port map(byteIn => t0_x1, byteOut => t0_x11);
    t1x11: x11 port map(byteIn => t1_x1, byteOut => t1_x11);
    t2x11: x11 port map(byteIn => t2_x1, byteOut => t2_x11);
    t3x11: x11 port map(byteIn => t3_x1, byteOut => t3_x11);

    t0x13: x13 port map(byteIn => t0_x1, byteOut => t0_x13);
    t1x13: x13 port map(byteIn => t1_x1, byteOut => t1_x13);
    t2x13: x13 port map(byteIn => t2_x1, byteOut => t2_x13);
    t3x13: x13 port map(byteIn => t3_x1, byteOut => t3_x13);
    
    t0x14: x14 port map(byteIn => t0_x1, byteOut => t0_x14);
    t1x14: x14 port map(byteIn => t1_x1, byteOut => t1_x14);
    t2x14: x14 port map(byteIn => t2_x1, byteOut => t2_x14);
    t3x14: x14 port map(byteIn => t3_x1, byteOut => t3_x14);

    wordOut(31 downto 24) <= t0_x14 XOR t1_x11 XOR t2_x13 XOR t3_x9;
    wordOut(23 downto 16) <= t0_x9  XOR t1_x14 XOR t2_x11 XOR t3_x13;
    wordOut(15 downto 8)  <= t0_x13 XOR t1_x9  XOR t2_x14 XOR t3_x11;
    wordOut(7 downto 0)   <= t0_x11 XOR t1_x13 XOR t2_x9  XOR t3_x14;

end Behavioral;
